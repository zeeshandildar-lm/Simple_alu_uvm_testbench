package simplealu_pkg;
    import uvm_pkg::*;
    `include "simplealu_sequencer.sv"
	`include "simplealu_monitor.sv"
	`include "simplealu_driver.sv"
	`include "simplealu_agent.sv"
	`include "simplealu_scoreboard.sv"
	`include "simplealu_config.sv"
	`include "simplealu_env.sv"
	`include "simplealu_test.sv"
endpackage