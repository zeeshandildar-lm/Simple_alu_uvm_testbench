class simplealu_configuration extends uvm_object;
	`uvm_object_utils(simplealu_configuration)

	function new(string name = "");
		super.new(name);
	endfunction: new
endclass: simplealu_configuration